module FA_dataflow (Cout, Sum,In1,In2,Cin);
input[31:0] In1,In2;
input Cin;
output Cout;
output[31:0] Sum;
assign {Cout,Sum}=In1+In2+Cin;
endmodule